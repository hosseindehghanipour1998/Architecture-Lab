`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:09:07 08/18/2020 
// Design Name: 
// Module Name:    Execute_Stage 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Execute_Stage(
	input [15:0] 	in_Read_Data_1,
	input [15:0] 	in_Read_Data_2,
	input [15:0] 	in_Immediate,
	input 		 	in_ALUSrc,
	input	[1:0]  	in_ALUOp,
	
	output [15:0]	O_ALUResult,
	output 			O_Zero,
    );


endmodule
