`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   19:01:26 08/25/2020
// Design Name:   MIPS
// Module Name:   G:/GitRepositories/8th Semester/Architecture Lab 2020/MIPS/Codes/MIPS_Test_2.v
// Project Name:  MIPS
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: MIPS
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module MIPS_Test_2;

	// Inputs
	reg clk;

	// Instantiate the Unit Under Test (UUT)
	MIPS uut (
		.clk(clk)
	);

	initial begin
		// Initialize Inputs
		clk = 0;


		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
always #10 clk = ~clk;    
endmodule

